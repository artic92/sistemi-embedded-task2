----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:    12:14:52 06/26/2017
-- Design Name:
-- Module Name:    complex_abs - Structural
-- Project Name:
-- Target Devices:
-- Tool versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity complex_abs is
	 Generic ( complex_width : natural := 32 );
    Port ( clock : in STD_LOGIC;
					 reset_n : in STD_LOGIC;
					 input_value : in  STD_LOGIC_VECTOR (complex_width-1 downto 0);
           abs_value : out  STD_LOGIC_VECTOR ((complex_width/2)-1 downto 0));
end complex_abs;

architecture Structural of complex_abs is

component moltiplicatore_booth
generic (
  n : natural := 4;
  m : natural := 4
);
port (
  A       : in  STD_LOGIC_VECTOR (n-1 downto 0);
  B       : in  STD_LOGIC_VECTOR (m-1 downto 0);
  enable  : in  STD_LOGIC;
  reset_n : in  STD_LOGIC;
  clock   : in  STD_LOGIC;
  done    : out STD_LOGIC;
  P       : out STD_LOGIC_VECTOR (n+m-1 downto 0)
);
end component moltiplicatore_booth;


component ripple_carry_adder
generic (
  n : natural := 4
);
port (
  A     : in  STD_LOGIC_VECTOR (n-1 downto 0);
  B     : in  STD_LOGIC_VECTOR (n-1 downto 0);
  c_in  : in  STD_LOGIC;
  c_out : out STD_LOGIC;
  ovfl  : out STD_LOGIC;
  S     : out STD_LOGIC_VECTOR (n-1 downto 0)
);
end component ripple_carry_adder;

component square_root
generic (
  n : natural := 8
);
port (
  clock   : in  STD_LOGIC;
  reset_n : in  STD_LOGIC;
  enable  : in  STD_LOGIC;
  D       : in  STD_LOGIC_VECTOR (n-1 downto 0);
  root    : out STD_LOGIC_VECTOR ((n/2)-1 downto 0);
  done    : out STD_LOGIC
);
end component square_root;

component parte_controllo_complex_abs
port (
  clock       : in  STD_LOGIC;
  reset_n     : in  STD_LOGIC;
  done_mul    : in  STD_LOGIC;
  done_sqrt   : in  STD_LOGIC;
	reset_n_all : out STD_LOGIC;
  enable_mul  : out STD_LOGIC;
  enable_sqrt : out STD_LOGIC
);
end component parte_controllo_complex_abs;

signal en_mul_sig, en_sqrt_sig : std_logic;
signal done_real_sig, done_imag_sig, done_mul_sig, done_sqrt_sig : std_logic;
signal add_ovfl_sig, reset_n_all_sig : std_logic;
signal power_real_sig, power_imag_sig, res_add_sig : std_logic_vector(complex_width-1 downto 0);

begin

done_mul_sig <= done_real_sig and done_imag_sig;

multiplier_real : moltiplicatore_booth
generic map (
  n => (complex_width)/2,
  m => (complex_width)/2
)
port map (
  A       => input_value((complex_width/2)-1 downto 0),
  B       => input_value((complex_width/2)-1 downto 0),
  enable  => en_mul_sig,
  reset_n => reset_n_all_sig,
  clock   => clock,
  done    => done_real_sig,
  P       => power_real_sig
);

multiplier_imag : moltiplicatore_booth
generic map (
  n => (complex_width)/2,
  m => (complex_width)/2
)
port map (
  A       => input_value(complex_width-1 downto complex_width/2),
  B       => input_value(complex_width-1 downto complex_width/2),
  enable  => en_mul_sig,
  reset_n => reset_n_all_sig,
  clock   => clock,
  done    => done_imag_sig,
  P       => power_imag_sig
);

mul_res_add : ripple_carry_adder
generic map (
  n => complex_width
)
port map (
  A     => power_real_sig,
  B     => power_imag_sig,
  c_in  => '0',
  c_out => open,
  ovfl  => add_ovfl_sig,
  S     => res_add_sig
);

square_add_res : square_root
generic map (
	n => complex_width
)
port map (
	clock   => clock,
	reset_n => reset_n_all_sig,
	enable  => en_sqrt_sig,
	D       => res_add_sig,
	root    => abs_value,
	done    => done_sqrt_sig
);

control_unit : parte_controllo_complex_abs
port map (
  clock       => clock,
  reset_n     => reset_n,
  done_mul    => done_mul_sig,
  done_sqrt   => done_sqrt_sig,
	reset_n_all => reset_n_all_sig,
  enable_mul  => en_mul_sig,
  enable_sqrt => en_sqrt_sig
);

end Structural;
